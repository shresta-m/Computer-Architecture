`include "lab1.v"

module top;

reg [31:0] a, b;
wire [31:0] out;

ieee_adder adder (a,b,out);

initial
begin
	a = 32'b01010101010101010101010101010101; b = 32'b01010101001010101010101010101010;
	#5 a= 32'b01010101010101010101010101010101;b=32'b01010101010101010101010101010101;
	#10 a = 32'b11010101011111111101010101010100 ; b= 32'b01010100111111111111111010101110 ;
	// //a=32'b01000001000111000000000000000000;b=32'b00111111000100000000000000000000;
	#15a=32'b00111111000100000000000000000000;b=32'b01000001000111000000000000000000;//9.75,0.5625
	// answer : 0 10000010 01001010000000000000000
	#20 a=32'b11000000110001100110011001100110;b=32'b11000000001000000000000000000000 ; //-6.2,-2.5
	//answer : 1 10000010 00010110011001100110011
	
	// #10 a=32'b01000000001000000000000000000000;b=32'b00000000000000000000000000000000;// +ve,0
	// //#15 a=32'b11000000000100000000000000000000;b=32'b01000001000111000000000000000000;
	// #15 a = 32'b1_10000000_11100000000000000000000;b = 32'b0_10000000_11000000000000000000000;	//-3.37,3.5
	// #20 a = 32'b0_11111111_00000000000000000000000;b = 32'b1_11111100_00000000000000000000000;//infinity case
		
	

end
initial 
begin
	$monitor($time,"\na =      %b %b %b,\nb =      %b %b %b,\noutput = %b %b %b",a[31],a[30:23],a[22:0],b[31],b[30:23],b[22:0],out[31],out[30:23],out[22:0]);
	// $dumpfile("32bit_fadder.vcd");
    //     	$dumpvars;
end
endmodule


